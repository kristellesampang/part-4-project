-- Nios_System_2A.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios_System_2A is
	port (
		button_pio_external_connection_export : in    std_logic_vector(1 downto 0)  := (others => '0'); -- button_pio_external_connection.export
		button_pio_irq_irq                    : out   std_logic;                                        --                 button_pio_irq.irq
		clocks_ref_clk_clk                    : in    std_logic                     := '0';             --                 clocks_ref_clk.clk
		clocks_ref_reset_reset                : in    std_logic                     := '0';             --               clocks_ref_reset.reset
		clocks_sdram_clk_clk                  : out   std_logic;                                        --               clocks_sdram_clk.clk
		led_pio_external_connection_export    : out   std_logic_vector(7 downto 0);                     --    led_pio_external_connection.export
		sdram_wire_addr                       : out   std_logic_vector(12 downto 0);                    --                     sdram_wire.addr
		sdram_wire_ba                         : out   std_logic_vector(1 downto 0);                     --                               .ba
		sdram_wire_cas_n                      : out   std_logic;                                        --                               .cas_n
		sdram_wire_cke                        : out   std_logic;                                        --                               .cke
		sdram_wire_cs_n                       : out   std_logic;                                        --                               .cs_n
		sdram_wire_dq                         : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
		sdram_wire_dqm                        : out   std_logic_vector(1 downto 0);                     --                               .dqm
		sdram_wire_ras_n                      : out   std_logic;                                        --                               .ras_n
		sdram_wire_we_n                       : out   std_logic                                         --                               .we_n
	);
end entity Nios_System_2A;

architecture rtl of Nios_System_2A is
	component Nios_System_2A_BUTTON_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Nios_System_2A_BUTTON_pio;

	component top_level_systolic_array is
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			avs_control_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_control_write      : in  std_logic                     := 'X';             -- write
			avs_control_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_control_read       : in  std_logic                     := 'X';             -- read
			avs_control_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			avm_data_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_data_read          : out std_logic;                                        -- read
			avm_data_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_data_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_weight_address     : out std_logic_vector(31 downto 0);                    -- address
			avm_weight_read        : out std_logic;                                        -- read
			avm_weight_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_weight_waitrequest : in  std_logic                     := 'X'              -- waitrequest
		);
	end component top_level_systolic_array;

	component Nios_System_2A_DATA_BRAM is
		port (
			address     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_System_2A_DATA_BRAM;

	component Nios_System_2A_LED_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Nios_System_2A_LED_pio;

	component Nios_System_2A_WEIGHT_BRAM is
		port (
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_System_2A_WEIGHT_BRAM;

	component Nios_System_2A_clocks is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Nios_System_2A_clocks;

	component Nios_System_2A_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Nios_System_2A_cpu;

	component Nios_System_2A_high_res_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_System_2A_high_res_timer;

	component Nios_System_2A_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Nios_System_2A_jtag_uart;

	component Nios_System_2A_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_System_2A_onchip_memory;

	component Nios_System_2A_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Nios_System_2A_sdram;

	component Nios_System_2A_mm_interconnect_0 is
		port (
			clocks_sys_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			CustomTopLevel_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CustomTopLevel_0_data_address                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CustomTopLevel_0_data_waitrequest                  : out std_logic;                                        -- waitrequest
			CustomTopLevel_0_data_read                         : in  std_logic                     := 'X';             -- read
			CustomTopLevel_0_data_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			DATA_BRAM_s2_address                               : out std_logic_vector(3 downto 0);                     -- address
			DATA_BRAM_s2_write                                 : out std_logic;                                        -- write
			DATA_BRAM_s2_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DATA_BRAM_s2_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			DATA_BRAM_s2_byteenable                            : out std_logic_vector(3 downto 0);                     -- byteenable
			DATA_BRAM_s2_chipselect                            : out std_logic;                                        -- chipselect
			DATA_BRAM_s2_clken                                 : out std_logic                                         -- clken
		);
	end component Nios_System_2A_mm_interconnect_0;

	component Nios_System_2A_mm_interconnect_1 is
		port (
			clocks_sys_clk_clk                      : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			BUTTON_pio_s1_address                   : out std_logic_vector(1 downto 0);                     -- address
			BUTTON_pio_s1_write                     : out std_logic;                                        -- write
			BUTTON_pio_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			BUTTON_pio_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			BUTTON_pio_s1_chipselect                : out std_logic;                                        -- chipselect
			cpu_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			CustomTopLevel_0_control_address        : out std_logic_vector(2 downto 0);                     -- address
			CustomTopLevel_0_control_write          : out std_logic;                                        -- write
			CustomTopLevel_0_control_read           : out std_logic;                                        -- read
			CustomTopLevel_0_control_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CustomTopLevel_0_control_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			DATA_BRAM_s1_address                    : out std_logic_vector(3 downto 0);                     -- address
			DATA_BRAM_s1_write                      : out std_logic;                                        -- write
			DATA_BRAM_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DATA_BRAM_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			DATA_BRAM_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			DATA_BRAM_s1_chipselect                 : out std_logic;                                        -- chipselect
			DATA_BRAM_s1_clken                      : out std_logic;                                        -- clken
			high_res_timer_s1_address               : out std_logic_vector(2 downto 0);                     -- address
			high_res_timer_s1_write                 : out std_logic;                                        -- write
			high_res_timer_s1_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			high_res_timer_s1_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			high_res_timer_s1_chipselect            : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			LED_pio_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			LED_pio_s1_write                        : out std_logic;                                        -- write
			LED_pio_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_pio_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			LED_pio_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory_s1_address                : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory_s1_write                  : out std_logic;                                        -- write
			onchip_memory_s1_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                  : out std_logic;                                        -- clken
			sdram_s1_address                        : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                          : out std_logic;                                        -- write
			sdram_s1_read                           : out std_logic;                                        -- read
			sdram_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                     : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                     : out std_logic;                                        -- chipselect
			WEIGHT_BRAM_s1_address                  : out std_logic_vector(1 downto 0);                     -- address
			WEIGHT_BRAM_s1_write                    : out std_logic;                                        -- write
			WEIGHT_BRAM_s1_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			WEIGHT_BRAM_s1_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			WEIGHT_BRAM_s1_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			WEIGHT_BRAM_s1_chipselect               : out std_logic;                                        -- chipselect
			WEIGHT_BRAM_s1_clken                    : out std_logic                                         -- clken
		);
	end component Nios_System_2A_mm_interconnect_1;

	component Nios_System_2A_mm_interconnect_2 is
		port (
			clocks_sys_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			CustomTopLevel_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CustomTopLevel_0_weight_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CustomTopLevel_0_weight_waitrequest                : out std_logic;                                        -- waitrequest
			CustomTopLevel_0_weight_read                       : in  std_logic                     := 'X';             -- read
			CustomTopLevel_0_weight_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			WEIGHT_BRAM_s2_address                             : out std_logic_vector(1 downto 0);                     -- address
			WEIGHT_BRAM_s2_write                               : out std_logic;                                        -- write
			WEIGHT_BRAM_s2_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			WEIGHT_BRAM_s2_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			WEIGHT_BRAM_s2_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			WEIGHT_BRAM_s2_chipselect                          : out std_logic;                                        -- chipselect
			WEIGHT_BRAM_s2_clken                               : out std_logic                                         -- clken
		);
	end component Nios_System_2A_mm_interconnect_2;

	component Nios_System_2A_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Nios_System_2A_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clocks_sys_clk_clk                                            : std_logic;                     -- clocks:sys_clk_clk -> [BUTTON_pio:clk, CustomTopLevel_0:clk, DATA_BRAM:clk, LED_pio:clk, WEIGHT_BRAM:clk, cpu:clk, high_res_timer:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:clocks_sys_clk_clk, mm_interconnect_1:clocks_sys_clk_clk, mm_interconnect_2:clocks_sys_clk_clk, onchip_memory:clk, rst_controller:clk, sdram:clk]
	signal customtoplevel_0_data_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:CustomTopLevel_0_data_readdata -> CustomTopLevel_0:avm_data_readdata
	signal customtoplevel_0_data_waitrequest                             : std_logic;                     -- mm_interconnect_0:CustomTopLevel_0_data_waitrequest -> CustomTopLevel_0:avm_data_waitrequest
	signal customtoplevel_0_data_address                                 : std_logic_vector(31 downto 0); -- CustomTopLevel_0:avm_data_address -> mm_interconnect_0:CustomTopLevel_0_data_address
	signal customtoplevel_0_data_read                                    : std_logic;                     -- CustomTopLevel_0:avm_data_read -> mm_interconnect_0:CustomTopLevel_0_data_read
	signal mm_interconnect_0_data_bram_s2_chipselect                     : std_logic;                     -- mm_interconnect_0:DATA_BRAM_s2_chipselect -> DATA_BRAM:chipselect2
	signal mm_interconnect_0_data_bram_s2_readdata                       : std_logic_vector(31 downto 0); -- DATA_BRAM:readdata2 -> mm_interconnect_0:DATA_BRAM_s2_readdata
	signal mm_interconnect_0_data_bram_s2_address                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:DATA_BRAM_s2_address -> DATA_BRAM:address2
	signal mm_interconnect_0_data_bram_s2_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:DATA_BRAM_s2_byteenable -> DATA_BRAM:byteenable2
	signal mm_interconnect_0_data_bram_s2_write                          : std_logic;                     -- mm_interconnect_0:DATA_BRAM_s2_write -> DATA_BRAM:write2
	signal mm_interconnect_0_data_bram_s2_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:DATA_BRAM_s2_writedata -> DATA_BRAM:writedata2
	signal mm_interconnect_0_data_bram_s2_clken                          : std_logic;                     -- mm_interconnect_0:DATA_BRAM_s2_clken -> DATA_BRAM:clken2
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_1:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_1:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_1:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_1:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_1:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_1:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_1:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_customtoplevel_0_control_readdata           : std_logic_vector(31 downto 0); -- CustomTopLevel_0:avs_control_readdata -> mm_interconnect_1:CustomTopLevel_0_control_readdata
	signal mm_interconnect_1_customtoplevel_0_control_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_1:CustomTopLevel_0_control_address -> CustomTopLevel_0:avs_control_address
	signal mm_interconnect_1_customtoplevel_0_control_read               : std_logic;                     -- mm_interconnect_1:CustomTopLevel_0_control_read -> CustomTopLevel_0:avs_control_read
	signal mm_interconnect_1_customtoplevel_0_control_write              : std_logic;                     -- mm_interconnect_1:CustomTopLevel_0_control_write -> CustomTopLevel_0:avs_control_write
	signal mm_interconnect_1_customtoplevel_0_control_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_1:CustomTopLevel_0_control_writedata -> CustomTopLevel_0:avs_control_writedata
	signal mm_interconnect_1_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_1:cpu_debug_mem_slave_readdata
	signal mm_interconnect_1_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_1:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_1_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_1:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_1_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_1:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_1_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_1:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_1_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_1:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_1_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_1:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_1_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_1_onchip_memory_s1_chipselect                 : std_logic;                     -- mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_1_onchip_memory_s1_readdata                   : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	signal mm_interconnect_1_onchip_memory_s1_address                    : std_logic_vector(12 downto 0); -- mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_1_onchip_memory_s1_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_1_onchip_memory_s1_write                      : std_logic;                     -- mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_1_onchip_memory_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_1_onchip_memory_s1_clken                      : std_logic;                     -- mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_1_high_res_timer_s1_chipselect                : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	signal mm_interconnect_1_high_res_timer_s1_readdata                  : std_logic_vector(15 downto 0); -- high_res_timer:readdata -> mm_interconnect_1:high_res_timer_s1_readdata
	signal mm_interconnect_1_high_res_timer_s1_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_1:high_res_timer_s1_address -> high_res_timer:address
	signal mm_interconnect_1_high_res_timer_s1_write                     : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_write -> mm_interconnect_1_high_res_timer_s1_write:in
	signal mm_interconnect_1_high_res_timer_s1_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_1:high_res_timer_s1_writedata -> high_res_timer:writedata
	signal mm_interconnect_1_button_pio_s1_chipselect                    : std_logic;                     -- mm_interconnect_1:BUTTON_pio_s1_chipselect -> BUTTON_pio:chipselect
	signal mm_interconnect_1_button_pio_s1_readdata                      : std_logic_vector(31 downto 0); -- BUTTON_pio:readdata -> mm_interconnect_1:BUTTON_pio_s1_readdata
	signal mm_interconnect_1_button_pio_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:BUTTON_pio_s1_address -> BUTTON_pio:address
	signal mm_interconnect_1_button_pio_s1_write                         : std_logic;                     -- mm_interconnect_1:BUTTON_pio_s1_write -> mm_interconnect_1_button_pio_s1_write:in
	signal mm_interconnect_1_button_pio_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_1:BUTTON_pio_s1_writedata -> BUTTON_pio:writedata
	signal mm_interconnect_1_led_pio_s1_chipselect                       : std_logic;                     -- mm_interconnect_1:LED_pio_s1_chipselect -> LED_pio:chipselect
	signal mm_interconnect_1_led_pio_s1_readdata                         : std_logic_vector(31 downto 0); -- LED_pio:readdata -> mm_interconnect_1:LED_pio_s1_readdata
	signal mm_interconnect_1_led_pio_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_1:LED_pio_s1_address -> LED_pio:address
	signal mm_interconnect_1_led_pio_s1_write                            : std_logic;                     -- mm_interconnect_1:LED_pio_s1_write -> mm_interconnect_1_led_pio_s1_write:in
	signal mm_interconnect_1_led_pio_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:LED_pio_s1_writedata -> LED_pio:writedata
	signal mm_interconnect_1_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_1_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	signal mm_interconnect_1_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	signal mm_interconnect_1_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_1_sdram_s1_read                               : std_logic;                     -- mm_interconnect_1:sdram_s1_read -> mm_interconnect_1_sdram_s1_read:in
	signal mm_interconnect_1_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sdram_s1_byteenable -> mm_interconnect_1_sdram_s1_byteenable:in
	signal mm_interconnect_1_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	signal mm_interconnect_1_sdram_s1_write                              : std_logic;                     -- mm_interconnect_1:sdram_s1_write -> mm_interconnect_1_sdram_s1_write:in
	signal mm_interconnect_1_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_1_data_bram_s1_chipselect                     : std_logic;                     -- mm_interconnect_1:DATA_BRAM_s1_chipselect -> DATA_BRAM:chipselect
	signal mm_interconnect_1_data_bram_s1_readdata                       : std_logic_vector(31 downto 0); -- DATA_BRAM:readdata -> mm_interconnect_1:DATA_BRAM_s1_readdata
	signal mm_interconnect_1_data_bram_s1_address                        : std_logic_vector(3 downto 0);  -- mm_interconnect_1:DATA_BRAM_s1_address -> DATA_BRAM:address
	signal mm_interconnect_1_data_bram_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_1:DATA_BRAM_s1_byteenable -> DATA_BRAM:byteenable
	signal mm_interconnect_1_data_bram_s1_write                          : std_logic;                     -- mm_interconnect_1:DATA_BRAM_s1_write -> DATA_BRAM:write
	signal mm_interconnect_1_data_bram_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:DATA_BRAM_s1_writedata -> DATA_BRAM:writedata
	signal mm_interconnect_1_data_bram_s1_clken                          : std_logic;                     -- mm_interconnect_1:DATA_BRAM_s1_clken -> DATA_BRAM:clken
	signal mm_interconnect_1_weight_bram_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:WEIGHT_BRAM_s1_chipselect -> WEIGHT_BRAM:chipselect
	signal mm_interconnect_1_weight_bram_s1_readdata                     : std_logic_vector(31 downto 0); -- WEIGHT_BRAM:readdata -> mm_interconnect_1:WEIGHT_BRAM_s1_readdata
	signal mm_interconnect_1_weight_bram_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:WEIGHT_BRAM_s1_address -> WEIGHT_BRAM:address
	signal mm_interconnect_1_weight_bram_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:WEIGHT_BRAM_s1_byteenable -> WEIGHT_BRAM:byteenable
	signal mm_interconnect_1_weight_bram_s1_write                        : std_logic;                     -- mm_interconnect_1:WEIGHT_BRAM_s1_write -> WEIGHT_BRAM:write
	signal mm_interconnect_1_weight_bram_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:WEIGHT_BRAM_s1_writedata -> WEIGHT_BRAM:writedata
	signal mm_interconnect_1_weight_bram_s1_clken                        : std_logic;                     -- mm_interconnect_1:WEIGHT_BRAM_s1_clken -> WEIGHT_BRAM:clken
	signal customtoplevel_0_weight_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_2:CustomTopLevel_0_weight_readdata -> CustomTopLevel_0:avm_weight_readdata
	signal customtoplevel_0_weight_waitrequest                           : std_logic;                     -- mm_interconnect_2:CustomTopLevel_0_weight_waitrequest -> CustomTopLevel_0:avm_weight_waitrequest
	signal customtoplevel_0_weight_address                               : std_logic_vector(31 downto 0); -- CustomTopLevel_0:avm_weight_address -> mm_interconnect_2:CustomTopLevel_0_weight_address
	signal customtoplevel_0_weight_read                                  : std_logic;                     -- CustomTopLevel_0:avm_weight_read -> mm_interconnect_2:CustomTopLevel_0_weight_read
	signal mm_interconnect_2_weight_bram_s2_chipselect                   : std_logic;                     -- mm_interconnect_2:WEIGHT_BRAM_s2_chipselect -> WEIGHT_BRAM:chipselect2
	signal mm_interconnect_2_weight_bram_s2_readdata                     : std_logic_vector(31 downto 0); -- WEIGHT_BRAM:readdata2 -> mm_interconnect_2:WEIGHT_BRAM_s2_readdata
	signal mm_interconnect_2_weight_bram_s2_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_2:WEIGHT_BRAM_s2_address -> WEIGHT_BRAM:address2
	signal mm_interconnect_2_weight_bram_s2_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_2:WEIGHT_BRAM_s2_byteenable -> WEIGHT_BRAM:byteenable2
	signal mm_interconnect_2_weight_bram_s2_write                        : std_logic;                     -- mm_interconnect_2:WEIGHT_BRAM_s2_write -> WEIGHT_BRAM:write2
	signal mm_interconnect_2_weight_bram_s2_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_2:WEIGHT_BRAM_s2_writedata -> WEIGHT_BRAM:writedata2
	signal mm_interconnect_2_weight_bram_s2_clken                        : std_logic;                     -- mm_interconnect_2:WEIGHT_BRAM_s2_clken -> WEIGHT_BRAM:clken2
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- high_res_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [CustomTopLevel_0:reset, DATA_BRAM:reset, WEIGHT_BRAM:reset, irq_mapper:reset, mm_interconnect_0:CustomTopLevel_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_2:CustomTopLevel_0_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [DATA_BRAM:reset_req, WEIGHT_BRAM:reset_req, cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                 : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in0
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_1_high_res_timer_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_1_high_res_timer_s1_write:inv -> high_res_timer:write_n
	signal mm_interconnect_1_button_pio_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_1_button_pio_s1_write:inv -> BUTTON_pio:write_n
	signal mm_interconnect_1_led_pio_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_1_led_pio_s1_write:inv -> LED_pio:write_n
	signal mm_interconnect_1_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_1_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_1_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_1_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_1_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_1_sdram_s1_write:inv -> sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [BUTTON_pio:reset_n, LED_pio:reset_n, cpu:reset_n, high_res_timer:reset_n, jtag_uart:rst_n, sdram:reset_n]

begin

	button_pio : component Nios_System_2A_BUTTON_pio
		port map (
			clk        => clocks_sys_clk_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_1_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_external_connection_export,           -- external_connection.export
			irq        => button_pio_irq_irq                               --                 irq.irq
		);

	customtoplevel_0 : component top_level_systolic_array
		port map (
			clk                    => clocks_sys_clk_clk,                                   --   clock.clk
			reset                  => rst_controller_reset_out_reset,                       --   reset.reset
			avs_control_address    => mm_interconnect_1_customtoplevel_0_control_address,   -- control.address
			avs_control_write      => mm_interconnect_1_customtoplevel_0_control_write,     --        .write
			avs_control_writedata  => mm_interconnect_1_customtoplevel_0_control_writedata, --        .writedata
			avs_control_read       => mm_interconnect_1_customtoplevel_0_control_read,      --        .read
			avs_control_readdata   => mm_interconnect_1_customtoplevel_0_control_readdata,  --        .readdata
			avm_data_address       => customtoplevel_0_data_address,                        --    data.address
			avm_data_read          => customtoplevel_0_data_read,                           --        .read
			avm_data_readdata      => customtoplevel_0_data_readdata,                       --        .readdata
			avm_data_waitrequest   => customtoplevel_0_data_waitrequest,                    --        .waitrequest
			avm_weight_address     => customtoplevel_0_weight_address,                      --  weight.address
			avm_weight_read        => customtoplevel_0_weight_read,                         --        .read
			avm_weight_readdata    => customtoplevel_0_weight_readdata,                     --        .readdata
			avm_weight_waitrequest => customtoplevel_0_weight_waitrequest                   --        .waitrequest
		);

	data_bram : component Nios_System_2A_DATA_BRAM
		port map (
			address     => mm_interconnect_1_data_bram_s1_address,    --     s1.address
			clken       => mm_interconnect_1_data_bram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_data_bram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_data_bram_s1_write,      --       .write
			readdata    => mm_interconnect_1_data_bram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_data_bram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_data_bram_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_0_data_bram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_data_bram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_data_bram_s2_clken,      --       .clken
			write2      => mm_interconnect_0_data_bram_s2_write,      --       .write
			readdata2   => mm_interconnect_0_data_bram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_data_bram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_data_bram_s2_byteenable, --       .byteenable
			clk         => clocks_sys_clk_clk,                        --   clk1.clk
			reset       => rst_controller_reset_out_reset,            -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,        --       .reset_req
			freeze      => '0'                                        -- (terminated)
		);

	led_pio : component Nios_System_2A_LED_pio
		port map (
			clk        => clocks_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	weight_bram : component Nios_System_2A_WEIGHT_BRAM
		port map (
			address     => mm_interconnect_1_weight_bram_s1_address,    --     s1.address
			clken       => mm_interconnect_1_weight_bram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_weight_bram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_weight_bram_s1_write,      --       .write
			readdata    => mm_interconnect_1_weight_bram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_weight_bram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_weight_bram_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_2_weight_bram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_2_weight_bram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_2_weight_bram_s2_clken,      --       .clken
			write2      => mm_interconnect_2_weight_bram_s2_write,      --       .write
			readdata2   => mm_interconnect_2_weight_bram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_2_weight_bram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_2_weight_bram_s2_byteenable, --       .byteenable
			clk         => clocks_sys_clk_clk,                          --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze      => '0'                                          -- (terminated)
		);

	clocks : component Nios_System_2A_clocks
		port map (
			ref_clk_clk        => clocks_ref_clk_clk,     --      ref_clk.clk
			ref_reset_reset    => clocks_ref_reset_reset, --    ref_reset.reset
			sys_clk_clk        => clocks_sys_clk_clk,     --      sys_clk.clk
			sdram_clk_clk      => clocks_sdram_clk_clk,   --    sdram_clk.clk
			reset_source_reset => open                    -- reset_source.reset
		);

	cpu : component Nios_System_2A_cpu
		port map (
			clk                                 => clocks_sys_clk_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	high_res_timer : component Nios_System_2A_high_res_timer
		port map (
			clk        => clocks_sys_clk_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_1_high_res_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_high_res_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_high_res_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_high_res_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_high_res_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                             --   irq.irq
		);

	jtag_uart : component Nios_System_2A_jtag_uart
		port map (
			clk            => clocks_sys_clk_clk,                                            --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	onchip_memory : component Nios_System_2A_onchip_memory
		port map (
			clk        => clocks_sys_clk_clk,                            --   clk1.clk
			address    => mm_interconnect_1_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_1_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_1_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	sdram : component Nios_System_2A_sdram
		port map (
			clk            => clocks_sys_clk_clk,                              --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_1_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_1_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_1_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_1_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_1_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_1_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_1_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_1_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_1_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	mm_interconnect_0 : component Nios_System_2A_mm_interconnect_0
		port map (
			clocks_sys_clk_clk                                 => clocks_sys_clk_clk,                        --                               clocks_sys_clk.clk
			CustomTopLevel_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,            -- CustomTopLevel_0_reset_reset_bridge_in_reset.reset
			CustomTopLevel_0_data_address                      => customtoplevel_0_data_address,             --                        CustomTopLevel_0_data.address
			CustomTopLevel_0_data_waitrequest                  => customtoplevel_0_data_waitrequest,         --                                             .waitrequest
			CustomTopLevel_0_data_read                         => customtoplevel_0_data_read,                --                                             .read
			CustomTopLevel_0_data_readdata                     => customtoplevel_0_data_readdata,            --                                             .readdata
			DATA_BRAM_s2_address                               => mm_interconnect_0_data_bram_s2_address,    --                                 DATA_BRAM_s2.address
			DATA_BRAM_s2_write                                 => mm_interconnect_0_data_bram_s2_write,      --                                             .write
			DATA_BRAM_s2_readdata                              => mm_interconnect_0_data_bram_s2_readdata,   --                                             .readdata
			DATA_BRAM_s2_writedata                             => mm_interconnect_0_data_bram_s2_writedata,  --                                             .writedata
			DATA_BRAM_s2_byteenable                            => mm_interconnect_0_data_bram_s2_byteenable, --                                             .byteenable
			DATA_BRAM_s2_chipselect                            => mm_interconnect_0_data_bram_s2_chipselect, --                                             .chipselect
			DATA_BRAM_s2_clken                                 => mm_interconnect_0_data_bram_s2_clken       --                                             .clken
		);

	mm_interconnect_1 : component Nios_System_2A_mm_interconnect_1
		port map (
			clocks_sys_clk_clk                      => clocks_sys_clk_clk,                                        --                  clocks_sys_clk.clk
			cpu_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            -- cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                                   --                 cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                                --                                .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                                      --                                .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                                  --                                .readdata
			cpu_data_master_readdatavalid           => cpu_data_master_readdatavalid,                             --                                .readdatavalid
			cpu_data_master_write                   => cpu_data_master_write,                                     --                                .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                                 --                                .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                            --          cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                               --                                .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                .readdata
			cpu_instruction_master_readdatavalid    => cpu_instruction_master_readdatavalid,                      --                                .readdatavalid
			BUTTON_pio_s1_address                   => mm_interconnect_1_button_pio_s1_address,                   --                   BUTTON_pio_s1.address
			BUTTON_pio_s1_write                     => mm_interconnect_1_button_pio_s1_write,                     --                                .write
			BUTTON_pio_s1_readdata                  => mm_interconnect_1_button_pio_s1_readdata,                  --                                .readdata
			BUTTON_pio_s1_writedata                 => mm_interconnect_1_button_pio_s1_writedata,                 --                                .writedata
			BUTTON_pio_s1_chipselect                => mm_interconnect_1_button_pio_s1_chipselect,                --                                .chipselect
			cpu_debug_mem_slave_address             => mm_interconnect_1_cpu_debug_mem_slave_address,             --             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write               => mm_interconnect_1_cpu_debug_mem_slave_write,               --                                .write
			cpu_debug_mem_slave_read                => mm_interconnect_1_cpu_debug_mem_slave_read,                --                                .read
			cpu_debug_mem_slave_readdata            => mm_interconnect_1_cpu_debug_mem_slave_readdata,            --                                .readdata
			cpu_debug_mem_slave_writedata           => mm_interconnect_1_cpu_debug_mem_slave_writedata,           --                                .writedata
			cpu_debug_mem_slave_byteenable          => mm_interconnect_1_cpu_debug_mem_slave_byteenable,          --                                .byteenable
			cpu_debug_mem_slave_waitrequest         => mm_interconnect_1_cpu_debug_mem_slave_waitrequest,         --                                .waitrequest
			cpu_debug_mem_slave_debugaccess         => mm_interconnect_1_cpu_debug_mem_slave_debugaccess,         --                                .debugaccess
			CustomTopLevel_0_control_address        => mm_interconnect_1_customtoplevel_0_control_address,        --        CustomTopLevel_0_control.address
			CustomTopLevel_0_control_write          => mm_interconnect_1_customtoplevel_0_control_write,          --                                .write
			CustomTopLevel_0_control_read           => mm_interconnect_1_customtoplevel_0_control_read,           --                                .read
			CustomTopLevel_0_control_readdata       => mm_interconnect_1_customtoplevel_0_control_readdata,       --                                .readdata
			CustomTopLevel_0_control_writedata      => mm_interconnect_1_customtoplevel_0_control_writedata,      --                                .writedata
			DATA_BRAM_s1_address                    => mm_interconnect_1_data_bram_s1_address,                    --                    DATA_BRAM_s1.address
			DATA_BRAM_s1_write                      => mm_interconnect_1_data_bram_s1_write,                      --                                .write
			DATA_BRAM_s1_readdata                   => mm_interconnect_1_data_bram_s1_readdata,                   --                                .readdata
			DATA_BRAM_s1_writedata                  => mm_interconnect_1_data_bram_s1_writedata,                  --                                .writedata
			DATA_BRAM_s1_byteenable                 => mm_interconnect_1_data_bram_s1_byteenable,                 --                                .byteenable
			DATA_BRAM_s1_chipselect                 => mm_interconnect_1_data_bram_s1_chipselect,                 --                                .chipselect
			DATA_BRAM_s1_clken                      => mm_interconnect_1_data_bram_s1_clken,                      --                                .clken
			high_res_timer_s1_address               => mm_interconnect_1_high_res_timer_s1_address,               --               high_res_timer_s1.address
			high_res_timer_s1_write                 => mm_interconnect_1_high_res_timer_s1_write,                 --                                .write
			high_res_timer_s1_readdata              => mm_interconnect_1_high_res_timer_s1_readdata,              --                                .readdata
			high_res_timer_s1_writedata             => mm_interconnect_1_high_res_timer_s1_writedata,             --                                .writedata
			high_res_timer_s1_chipselect            => mm_interconnect_1_high_res_timer_s1_chipselect,            --                                .chipselect
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,     --     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,       --                                .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,        --                                .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,  --                                .chipselect
			LED_pio_s1_address                      => mm_interconnect_1_led_pio_s1_address,                      --                      LED_pio_s1.address
			LED_pio_s1_write                        => mm_interconnect_1_led_pio_s1_write,                        --                                .write
			LED_pio_s1_readdata                     => mm_interconnect_1_led_pio_s1_readdata,                     --                                .readdata
			LED_pio_s1_writedata                    => mm_interconnect_1_led_pio_s1_writedata,                    --                                .writedata
			LED_pio_s1_chipselect                   => mm_interconnect_1_led_pio_s1_chipselect,                   --                                .chipselect
			onchip_memory_s1_address                => mm_interconnect_1_onchip_memory_s1_address,                --                onchip_memory_s1.address
			onchip_memory_s1_write                  => mm_interconnect_1_onchip_memory_s1_write,                  --                                .write
			onchip_memory_s1_readdata               => mm_interconnect_1_onchip_memory_s1_readdata,               --                                .readdata
			onchip_memory_s1_writedata              => mm_interconnect_1_onchip_memory_s1_writedata,              --                                .writedata
			onchip_memory_s1_byteenable             => mm_interconnect_1_onchip_memory_s1_byteenable,             --                                .byteenable
			onchip_memory_s1_chipselect             => mm_interconnect_1_onchip_memory_s1_chipselect,             --                                .chipselect
			onchip_memory_s1_clken                  => mm_interconnect_1_onchip_memory_s1_clken,                  --                                .clken
			sdram_s1_address                        => mm_interconnect_1_sdram_s1_address,                        --                        sdram_s1.address
			sdram_s1_write                          => mm_interconnect_1_sdram_s1_write,                          --                                .write
			sdram_s1_read                           => mm_interconnect_1_sdram_s1_read,                           --                                .read
			sdram_s1_readdata                       => mm_interconnect_1_sdram_s1_readdata,                       --                                .readdata
			sdram_s1_writedata                      => mm_interconnect_1_sdram_s1_writedata,                      --                                .writedata
			sdram_s1_byteenable                     => mm_interconnect_1_sdram_s1_byteenable,                     --                                .byteenable
			sdram_s1_readdatavalid                  => mm_interconnect_1_sdram_s1_readdatavalid,                  --                                .readdatavalid
			sdram_s1_waitrequest                    => mm_interconnect_1_sdram_s1_waitrequest,                    --                                .waitrequest
			sdram_s1_chipselect                     => mm_interconnect_1_sdram_s1_chipselect,                     --                                .chipselect
			WEIGHT_BRAM_s1_address                  => mm_interconnect_1_weight_bram_s1_address,                  --                  WEIGHT_BRAM_s1.address
			WEIGHT_BRAM_s1_write                    => mm_interconnect_1_weight_bram_s1_write,                    --                                .write
			WEIGHT_BRAM_s1_readdata                 => mm_interconnect_1_weight_bram_s1_readdata,                 --                                .readdata
			WEIGHT_BRAM_s1_writedata                => mm_interconnect_1_weight_bram_s1_writedata,                --                                .writedata
			WEIGHT_BRAM_s1_byteenable               => mm_interconnect_1_weight_bram_s1_byteenable,               --                                .byteenable
			WEIGHT_BRAM_s1_chipselect               => mm_interconnect_1_weight_bram_s1_chipselect,               --                                .chipselect
			WEIGHT_BRAM_s1_clken                    => mm_interconnect_1_weight_bram_s1_clken                     --                                .clken
		);

	mm_interconnect_2 : component Nios_System_2A_mm_interconnect_2
		port map (
			clocks_sys_clk_clk                                 => clocks_sys_clk_clk,                          --                               clocks_sys_clk.clk
			CustomTopLevel_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,              -- CustomTopLevel_0_reset_reset_bridge_in_reset.reset
			CustomTopLevel_0_weight_address                    => customtoplevel_0_weight_address,             --                      CustomTopLevel_0_weight.address
			CustomTopLevel_0_weight_waitrequest                => customtoplevel_0_weight_waitrequest,         --                                             .waitrequest
			CustomTopLevel_0_weight_read                       => customtoplevel_0_weight_read,                --                                             .read
			CustomTopLevel_0_weight_readdata                   => customtoplevel_0_weight_readdata,            --                                             .readdata
			WEIGHT_BRAM_s2_address                             => mm_interconnect_2_weight_bram_s2_address,    --                               WEIGHT_BRAM_s2.address
			WEIGHT_BRAM_s2_write                               => mm_interconnect_2_weight_bram_s2_write,      --                                             .write
			WEIGHT_BRAM_s2_readdata                            => mm_interconnect_2_weight_bram_s2_readdata,   --                                             .readdata
			WEIGHT_BRAM_s2_writedata                           => mm_interconnect_2_weight_bram_s2_writedata,  --                                             .writedata
			WEIGHT_BRAM_s2_byteenable                          => mm_interconnect_2_weight_bram_s2_byteenable, --                                             .byteenable
			WEIGHT_BRAM_s2_chipselect                          => mm_interconnect_2_weight_bram_s2_chipselect, --                                             .chipselect
			WEIGHT_BRAM_s2_clken                               => mm_interconnect_2_weight_bram_s2_clken       --                                             .clken
		);

	irq_mapper : component Nios_System_2A_irq_mapper
		port map (
			clk           => clocks_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,      -- reset_in0.reset
			clk            => clocks_sys_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_1_high_res_timer_s1_write_ports_inv <= not mm_interconnect_1_high_res_timer_s1_write;

	mm_interconnect_1_button_pio_s1_write_ports_inv <= not mm_interconnect_1_button_pio_s1_write;

	mm_interconnect_1_led_pio_s1_write_ports_inv <= not mm_interconnect_1_led_pio_s1_write;

	mm_interconnect_1_sdram_s1_read_ports_inv <= not mm_interconnect_1_sdram_s1_read;

	mm_interconnect_1_sdram_s1_byteenable_ports_inv <= not mm_interconnect_1_sdram_s1_byteenable;

	mm_interconnect_1_sdram_s1_write_ports_inv <= not mm_interconnect_1_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Nios_System_2A
